module mytext

pub fn hello() int {
	println('hello world')
	return 1
}
